class env_cfg_class;
bit [2:0] phase;
OS_type o_sets; 
GEN gen_speed;
tr_type transaction_type;
bit  data_income;  
endclass: env_cfg_class

