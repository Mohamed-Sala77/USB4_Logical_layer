package tb_pkg;
	

	// Transactions
	`include "elec_layer_tr.svh"
	`include "upper_layer_tr.svh"
	`include "config_space_pkg.sv"

	// Symbol Generator
	`include "symbols.svh"

	// Timing Parameters 
	`include "timing_parameters.svh"

	// REFERENCE MODEL
	`include "int_packet.sv"
	`include "R_Mod_extentions.sv"
	`include "my_memory.sv"
	`include "primary_steps.sv"

	`include "phase1.sv"
	`include "phase2.sv"
	`include "phase3.sv"
	`include "phase4.sv"
	`include "phase5.sv"

	`include "ref_model.sv"


	
	// Generators
	`include "upper_layer_generator.svh"
	`include "elec_layer_generator.svh"
	`include "config_space_stimulus_generator_pkg.sv"
	
	// Virtual Sequence
	`include "virtual_sequence_pkg.sv"

	// UPPER LAYER FILES
	`include "upper_layer_scoreboard.svh"
	`include "upper_layer_driver.svh"
	`include "upper_layer_monitor.svh"
	`include "upper_layer_agent.svh"


	// ELECTRICAL LAYER FILES	
	`include "elec_layer_driver.svh"
	`include "elec_layer_monitor.svh"
	`include "elec_layer_scoreboard.svh"
	`include "elec_layer_agent.svh"


	// CONFIGURATION SPACE LAYER FILES
	`include "config_space_driver_pkg.sv"
	`include "config_space_monitor_pkg.sv"
	`include "config_space_scoreboard_pkg.sv"
	`include "config_space_agent_pkg.sv"

	// ENVIRONMENT FILE
	`include "Environment.svh"
	
	// TEST FILE
	`include "Test.svh"




endpackage
