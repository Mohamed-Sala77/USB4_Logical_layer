///////////////////////****monitor package****//////////////////////////////
package electrical_layer_monitor_pkg;

	import electrical_layer_transaction_pkg::*;
	class electrical_layer_generator;
		// Declare your class variables, methods here
		
		 task run();
		 endtask
	endclass : electrical_layer_generator
	// Declare your data types, parameters, functions, tasks here
endpackage : electrical_layer_monitor_pkg