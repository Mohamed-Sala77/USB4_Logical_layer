
class mem;
bit   gen2 ;
bit   gen3 ;
bit   gen4 ;
bit [2:0]   gen_config ;
bit usb4;  // represent  the type of data that i should send to the scoreboard
                                    // 1 - it is  USB4 connection -/ 0- it is not USB4 connection
//bit [2:0] phase ;                  // represent the phase of the transaction

endclass //mem
