	parameter start_bit = 1'b0;
	parameter stop_bit = 1'b1;

	parameter [7:0] DLE = 8'hFE;	//Data Link Escape (DLE) Symbol – indicates the beginning of a Transaction. 
	parameter [7:0] ETX = 8'h40;	//End of Transaction (ETX) Symbol 

	parameter [7:0] LSE_lane0 = 8'b10000000;	//Lane State Event (LSE) - indicating LT_Fall for lane 0.
	parameter [7:0] LSE_lane1 = 8'b10100000;	//Lane State Event (LSE) - indicating LT_Fall for lane 1.

	parameter [7:0] STX_cmd = 8'b00000101;		//Start Transaction (STX) Symbol – defines the operation of the Transaction. 
	parameter [7:0] STX_rsp = 8'b00000100;		//Start Transaction (STX) Symbol – defines the operation of the Transaction. 


	//Constants sizes
	parameter TR_HEADER_SIZE = 20; 	// We need the first 20 bits of the transaction received to know the transaction type
	parameter MIN_TR_SIZE = 30;		//The minimum size of any transaction is 30 bits (LT Fall)
	parameter LT_TR_SIZE = 30;		//Size of the LT Transactions (30 bits)

	parameter SLOS_SIZE = 2112; // 66 * 32 = 2112 or 132 * 16 = 2112
	parameter TS_GEN_2_3_SIZE = 64;
	parameter TS_GEN_4_HEADER_SIZE = 28;
	parameter TS16_SIZE = 7168; // Size of 16 back to back TS (448 * 16 = 7168)

	parameter PRBS11_SYMBOL_SIZE = 420; // Size of the PRBS11 symbol
	parameter PRTS7_SYMBOL_SIZE = 420; // Size of the PRTS7 symbol




	//Ordered sets
	parameter [65:0] SLOS1_64 [31:0] = {66'b100100000000101000000100010000101010100100000001101000001110010001,
										66'b101011101011101010001010000101000100100010101101010000110000100111,
										66'b101001011100111001011110111001001010111011000010101110010000101110,
										66'b101001001010011011000111101110110010101011110000001001100001011111,
										66'b100010010001110110101101011000110001110111101101010010110000110011,
										66'b101001111110111100001010011001000111111010110000100011100101011011,
										66'b101000011010110011100011111011011000101101110100110101001111000011,
										66'b101001100110111111111010000000100100000101101000100110010101111110,
										66'b100001000011001010011111000111000110110110111011011010101101100000,
										66'b101101110001110101101101000110110010111011110010101001110000011101,
										66'b101000110101110111000101010110100000011001000011111010011000100111,
										66'b101101011100010001011010101001100000011111000011000110011110111111,
										66'b100010100001110001001101101011110110001001011101011001010001111000,
										66'b101011001101001111110011100001111011001100101111111100100000011101,
										66'b100000110100100111001101110111110101010001000000101010000100000100,
										66'b101010001011000101001110100011101001011010011001100111111111110000,
										66'b100000011000000011110000011001100011111111011000000101110000100101,
										66'b101001011001111001111100111100011110011011001111101111100010100011,
										66'b100100010111001010010111000110010110111110011010001111100101100011,
										66'b101001110110111101011010010001100110101111111000100000110101000111,
										66'b100000101101100100110111101111010010100100110001101111101110100010,
										66'b101010010100000110001000111101010110010000011110100011001001011111,
										66'b100110010001011110101001001000011011010011101100111010111110100010,
										66'b100010010101010110000000011100000011011000011101110011010101111100,
										66'b100001000110001010111101000010010010010110110110011011011111101101,
										66'b100000101100100100111101101110010110101110011000101111110100100001,
										66'b100011010010111100110010011111110111000001010110001000011101010011,
										66'b100100001111001001100111011111110101000001000010001010010101000110,
										66'b100000101111000100100110101101111000110100110111001111010111100100,
										66'b100100111010101110100000101001000100011010101011100000001011000001,
										66'b100011100010111011010010101100110000111111100110000011111100011000,
										66'b100110111100111010011110100111001001110111011101010101010000000000};


	parameter [2111:0] SLOS1_64_1 = {	SLOS1_64[0], SLOS1_64[1], SLOS1_64[2], SLOS1_64[3], SLOS1_64[4], SLOS1_64[5], SLOS1_64[6], SLOS1_64[7], 
										SLOS1_64[8], SLOS1_64[9], SLOS1_64[10], SLOS1_64[11], SLOS1_64[12], SLOS1_64[13], SLOS1_64[14], SLOS1_64[15], 
										SLOS1_64[16], SLOS1_64[17], SLOS1_64[18], SLOS1_64[19], SLOS1_64[20], SLOS1_64[21], SLOS1_64[22], SLOS1_64[23], 
										SLOS1_64[24], SLOS1_64[25], SLOS1_64[26], SLOS1_64[27], SLOS1_64[28], SLOS1_64[29], SLOS1_64[30], SLOS1_64[31]};


	parameter [65:0] SLOS2_64 [31:0] = {66'b101011111111010111111011101111010101011011111110010111110001101110,
										66'b100100010100010101110101111010111011011101010010101111001111011000,
										66'b100110100011000110100001000110110101000100111101010001101111010001,
										66'b100110110101100100111000010001001101010100001111110110011110100000,
										66'b101101101110001001010010100111001110001000010010101101001111001100,
										66'b100110000001000011110101100110111000000101001111011100011010100100,
										66'b100111100101001100011100000100100111010010001011001010110000111100,
										66'b100110011001000000000101111111011011111010010111011001101010000001,
										66'b101110111100110101100000111000111001001001000100100101010010011111,
										66'b100010001110001010010010111001001101000100001101010110001111100010,
										66'b100111001010001000111010101001011111100110111100000101100111011000,
										66'b100010100011101110100101010110011111100000111100111001100001000000,
										66'b101101011110001110110010010100001001110110100010100110101110000111,
										66'b100100110010110000001100011110000100110011010000000011011111100010,
										66'b101111001011011000110010001000001010101110111111010101111011111011,
										66'b100101110100111010110001011100010110100101100110011000000000001111,
										66'b101111100111111100001111100110011100000000100111111010001111011010,
										66'b100110100110000110000011000011100001100100110000010000011101011100,
										66'b101011101000110101101000111001101001000001100101110000011010011100,
										66'b100110001001000010100101101110011001010000000111011111001010111000,
										66'b101111010010011011001000010000101101011011001110010000010001011101,
										66'b100101101011111001110111000010101001101111100001011100110110100000,
										66'b101001101110100001010110110111100100101100010011000101000001011101,
										66'b101101101010101001111111100011111100100111100010001100101010000011,
										66'b101110111001110101000010111101101101101001001001100100100000010010,
										66'b101111010011011011000010010001101001010001100111010000001011011110,
										66'b101100101101000011001101100000001000111110101001110111100010101100,
										66'b101011110000110110011000100000001010111110111101110101101010111001,
										66'b101111010000111011011001010010000111001011001000110000101000011011,
										66'b101011000101010001011111010110111011100101010100011111110100111110,
										66'b101100011101000100101101010011001111000000011001111100000011100111,
										66'b101001000011000101100001011000110110001000100010101010101111111111};


	parameter [2111:0] SLOS2_64_1 = {	SLOS2_64[0], SLOS2_64[1], SLOS2_64[2], SLOS2_64[3], SLOS2_64[4], SLOS2_64[5], SLOS2_64[6], SLOS2_64[7], 
										SLOS2_64[8], SLOS2_64[9], SLOS2_64[10], SLOS2_64[11], SLOS2_64[12], SLOS2_64[13], SLOS2_64[14], SLOS2_64[15], 
										SLOS2_64[16], SLOS2_64[17], SLOS2_64[18], SLOS2_64[19], SLOS2_64[20], SLOS2_64[21], SLOS2_64[22], SLOS2_64[23], 
										SLOS2_64[24], SLOS2_64[25], SLOS2_64[26], SLOS2_64[27], SLOS2_64[28], SLOS2_64[29], SLOS2_64[30], SLOS2_64[31]};

	
	parameter [131:0] SLOS1_128 [15:0] = {	132'b101001000000001010000001000100001010101001000000011010000011100100011011101011101010001010000101000100100010101101010000110000100111,
											132'b101010010111001110010111101110010010101110110000101011100100001011101001001010011011000111101110110010101011110000001001100001011111,
											132'b101000100100011101101011010110001100011101111011010100101100001100111001111110111100001010011001000111111010110000100011100101011011,
											132'b101010000110101100111000111110110110001011011101001101010011110000111001100110111111111010000000100100000101101000100110010101111110,
											132'b101000010000110010100111110001110001101101101110110110101011011000001101110001110101101101000110110010111011110010101001110000011101,
											132'b101010001101011101110001010101101000000110010000111110100110001001111101011100010001011010101001100000011111000011000110011110111111,
											132'b101000101000011100010011011010111101100010010111010110010100011110001011001101001111110011100001111011001100101111111100100000011101,
											132'b101000001101001001110011011101111101010100010000001010100001000001001010001011000101001110100011101001011010011001100111111111110000,
											132'b101000000110000000111100000110011000111111110110000001011100001001011001011001111001111100111100011110011011001111101111100010100011,
											132'b101001000101110010100101110001100101101111100110100011111001011000111001110110111101011010010001100110101111111000100000110101000111,
											132'b101000001011011001001101111011110100101001001100011011111011101000101010010100000110001000111101010110010000011110100011001001011111,
											132'b101001100100010111101010010010000110110100111011001110101111101000100010010101010110000000011100000011011000011101110011010101111100,
											132'b101000010001100010101111010000100100100101101101100110110111111011010000101100100100111101101110010110101110011000101111110100100001,
											132'b101000110100101111001100100111111101110000010101100010000111010100110100001111001001100111011111110101000001000010001010010101000110,
											132'b101000001011110001001001101011011110001101001101110011110101111001000100111010101110100000101001000100011010101011100000001011000001,
											132'b101000111000101110110100101011001100001111111001100000111111000110000110111100111010011110100111001001110111011101010101010000000000};


	parameter [2111:0] SLOS1_128_1 = {	SLOS1_128[0], SLOS1_128[1], SLOS1_128[2], SLOS1_128[3], SLOS1_128[4], SLOS1_128[5], SLOS1_128[6], SLOS1_128[7], 
										SLOS1_128[8], SLOS1_128[9], SLOS1_128[10], SLOS1_128[11], SLOS1_128[12], SLOS1_128[13], SLOS1_128[14], SLOS1_128[15] };


	parameter [131:0] SLOS2_128 [15:0] = {	132'b101010111111110101111110111011110101010110111111100101111100011011100100010100010101110101111010111011011101010010101111001111011000,
											132'b101001101000110001101000010001101101010001001111010100011011110100010110110101100100111000010001001101010100001111110110011110100000,
											132'b101011011011100010010100101001110011100010000100101011010011110011000110000001000011110101100110111000000101001111011100011010100100,
											132'b101001111001010011000111000001001001110100100010110010101100001111000110011001000000000101111111011011111010010111011001101010000001,
											132'b101011101111001101011000001110001110010010010001001001010100100111110010001110001010010010111001001101000100001101010110001111100010,
											132'b101001110010100010001110101010010111111001101111000001011001110110000010100011101110100101010110011111100000111100111001100001000000,
											132'b101011010111100011101100100101000010011101101000101001101011100001110100110010110000001100011110000100110011010000000011011111100010,
											132'b101011110010110110001100100010000010101011101111110101011110111110110101110100111010110001011100010110100101100110011000000000001111,
											132'b101011111001111111000011111001100111000000001001111110100011110110100110100110000110000011000011100001100100110000010000011101011100,
											132'b101010111010001101011010001110011010010000011001011100000110100111000110001001000010100101101110011001010000000111011111001010111000,
											132'b101011110100100110110010000100001011010110110011100100000100010111010101101011111001110111000010101001101111100001011100110110100000,
											132'b101010011011101000010101101101111001001011000100110001010000010111011101101010101001111111100011111100100111100010001100101010000011,
											132'b101011101110011101010000101111011011011010010010011001001000000100101111010011011011000010010001101001010001100111010000001011011110,
											132'b101011001011010000110011011000000010001111101010011101111000101011001011110000110110011000100000001010111110111101110101101010111001,
											132'b101011110100001110110110010100100001110010110010001100001010000110111011000101010001011111010110111011100101010100011111110100111110,
											132'b101011000111010001001011010100110011110000000110011111000000111001111001000011000101100001011000110110001000100010101010101111111111};


	parameter [2111:0] SLOS2_128_1 = {	SLOS2_128[0], SLOS2_128[1], SLOS2_128[2], SLOS2_128[3], SLOS2_128[4], SLOS2_128[5], SLOS2_128[6], SLOS2_128[7], 
										SLOS2_128[8], SLOS2_128[9], SLOS2_128[10], SLOS2_128[11], SLOS2_128[12], SLOS2_128[13], SLOS2_128[14], SLOS2_128[15] };


	//Parameters for TS1 and TS2 symbols for Gen 2 and Gen 3
	parameter [7:0] lane_number_0 = 8'h00, lane_number_1 = 8'h01; // To indicate the lane number (one for lane 0  and one for lane 1)
	parameter [5:0] TSID_TS1 = 6'b100110; // To indicate TS1
	parameter [5:0] TSID_TS2 = 6'b011001; // To indicate TS2
	parameter [9:0] SCR = 10'b0011110010;

	//Parameters for TS symbols for Gen 4
	parameter [11:0] CURSOR = 12'h7E0;


	// Seeds for the Pseudo Random Sequences
	parameter [10:0] PRBS11_lane0_seed = 11'b11111111111;
	parameter [10:0] PRBS11_lane1_seed = 11'b11101110000;

	parameter [13:0] PRTS7_lane0_seed = 14'b01010101010101;
	parameter [13:0] PRTS7_lane1_seed = 14'b00_01_10_00_10_01_00;


	class TS_Symbols;
		
		bit TS1_lane_0_16 [$];
		bit TS1_lane_1_16 [$];
		bit [0:1] TS_234_lane_0_16 [$];
		bit [1:0] TS_234_lane_1_16 [$];

		bit [419:0] TS1_lane_0 [15:0];
		bit [419:0] TS1_lane_1 [15:0];
		bit [419:0] TS_234_lane_0 [15:0];
		bit [419:0] TS_234_lane_1 [15:0];

		

		task calculate_TS;

			int index = 28; 
			int indextrit = 28;
			
			PRBS11(TS16_SIZE, PRBS11_lane0_seed, TS1_lane_0_16);
			PRBS11(TS16_SIZE, PRBS11_lane1_seed, TS1_lane_1_16);
			PRTS7(TS16_SIZE/2, PRTS7_lane0_seed, TS_234_lane_0_16);
			PRTS7(TS16_SIZE/2, PRTS7_lane1_seed, TS_234_lane_1_16);
		

			for (int i = 0 ; i < 15; i++ )
			begin
				TS1_lane_0 [i] = { >> {TS1_lane_0_16 [index:index+419]} };
				TS1_lane_1 [i] = { >> {TS1_lane_1_16 [index:index+419]} };
				TS_234_lane_0 [i] = { >> {TS_234_lane_0_16 [indextrit:indextrit+209]} };
				TS_234_lane_1 [i] = { >> {TS_234_lane_1_16 [indextrit:indextrit+209]} };

				index += 419 + 29;
				indextrit += 209 + 15; // check numbers 209 & 15

			end

			// TS_234_lane_0[10] = TS_234_lane_0[0];
			// TS_234_lane_0[0] = 0;

			// TS_234_lane_1[10] = TS_234_lane_1[0];
			// TS_234_lane_1[0] = 0;

			// TS1_lane_0[10] = TS1_lane_0[0];
			// TS1_lane_0[0] = 0;

			//$display("TASK: TS2_Lane0 complete: %p",TS_234_lane_0_16);
			//$display("TASK: TS2_Lane1 complete: %p",TS_234_lane_1_16);
			//$display("TASK: TS1_Lane0: %b",TS1_lane_0 [0]);
			//$display("TASK: TS1_Lane1: %b",TS1_lane_1 [0]);

			//$display("[SYMBOLS] TASK: TS2_Lane0: %b",TS_234_lane_0 [0]);
			//$display("[SYMBOLS] TASK: TS2_Lane1: %b",TS_234_lane_1 [0]);
			
			//$stop;

		endtask

	endclass : TS_Symbols

	task PRBS11 (input int size ,input bit [10:0] seed, output bit PRBS11_INTERNAL [$]);

			//bit PRBS11_INTERNAL [$];
			bit [10:0] internal_reg;
			bit internal_bit10; bit internal_bit8;
			
			// repeat(size)
			// begin
			// 	void'(PRBS11_INTERNAL.pop_front());
			// end

			PRBS11_INTERNAL = {};

			internal_reg = seed;

			while (PRBS11_INTERNAL.size() != size)
			begin


				PRBS11_INTERNAL.push_back(internal_reg[10]);
				internal_bit8 = internal_reg[8]; 
				internal_bit10 = internal_reg[10];

				internal_reg[10] = internal_reg[9];
				internal_reg[9] = internal_reg[8];
				internal_reg[8] = internal_reg[7];
				internal_reg[7] = internal_reg[6];
				internal_reg[6] = internal_reg[5];
				internal_reg[5] = internal_reg[4];
				internal_reg[4] = internal_reg[3];
				internal_reg[3] = internal_reg[2];
				internal_reg[2] = internal_reg[1];
				internal_reg[1] = internal_reg[0];
				internal_reg[0] =  internal_bit8 ^ internal_bit10;

			end



			//$display("************************************************************");
			//$display("PRBS_INTERNAL11 : [%0p]",PRBS11_INTERNAL);
			//$display("************************************************************");


		endtask

		function bit[1:0] GF3 (input [1:0] A, input string op,input [1:0] B);
			case (op)
				"+":
				begin
					case({A,B})
						4'b00_00, 4'b01_10 , 4'b10_01:
						begin
							GF3 = 2'b00;
						end

						4'b00_01, 4'b01_00, 4'b10_10:
						begin
							GF3 = 2'b01;
						end

						4'b00_10, 4'b10_00, 4'b01_01:
						begin
							GF3 = 2'b10;
						end
					endcase
				end

				"*":
				begin
					case({A,B})
						4'b00_00 ,4'b00_01, 4'b00_10, 4'b01_00, 4'b10_00:
						begin
							GF3 = 2'b00;
						end

						4'b01_01, 4'b10_10:
						begin
							GF3 = 2'b01;
						end

						4'b10_01, 4'b01_10:
						begin
							GF3 = 2'b10;
						end
					endcase
				end

			endcase
		endfunction : GF3


		task PRTS7 (input int size, input bit[13:0] seed, output bit[1:0] PRBS7_INTERNAL [$] );

			//bit [1:0] PRBS7_INTERNAL [$];
			bit [13:0] internal_reg;
			bit [1:0] internal_trit2; bit[1:0] internal_trit7;
			// repeat(size)
			// begin
			// 	void'(PRBS7_INTERNAL.pop_front());
			// end

			PRBS7_INTERNAL = {};
			//$display("PRBS7_INTERNAL [%p]",PRBS7_INTERNAL);
			internal_reg = seed;
			while (PRBS7_INTERNAL.size() != size)
			begin


				PRBS7_INTERNAL.push_back(internal_reg[13:12]);
				internal_trit2 = internal_reg[3:2]; 
				internal_trit7 = GF3(2'b10,"*",internal_reg[13:12]);


				internal_reg[13:12] = internal_reg[11:10];
				internal_reg[11:10] = internal_reg[9:8];
				internal_reg[9:8] = internal_reg[7:6];
				internal_reg[7:6] = internal_reg[5:4];
				internal_reg[5:4] = internal_reg[3:2];
				internal_reg[3:2] = internal_reg[1:0];
				
				internal_reg[1:0] =  GF3( internal_trit2,"+", internal_trit7);

			end

			//$display("PRBS7_INTERNAL : [%0p]",PRBS7_INTERNAL);

		endtask

